//freq_show.v

module freq_show(
freq,

);
input [9:0]	freq;

//-----------------------------------

wire [3:0] 

endmodule
